`timescale 1ns / 1ps
module testbench_CheckParity(
    );

	reg [1:12] dataIn;
	wire [1:8] dataOut;
	integer result=0;
	//instances
	CheckParity ins( dataIn,   dataOut);	
	

	initial begin
	$display("Starting Testbench");
	
	#1;
	dataIn=12'b110000010100;
	#1;
	if (dataOut==8'b00000100) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00000100);
	#1;
	dataIn=12'b110100001001;
	#1;
	if (dataOut==8'b00001001) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00001001);
	#1;
	dataIn=12'b011100100110;
	#1;
	if (dataOut==8'b00010110) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00010110);
	#1;
	dataIn=12'b100100111011;
	#1;
	if (dataOut==8'b00011011) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00011011);
	#1;
	dataIn=12'b000111010100;
	#1;
	if (dataOut==8'b00100100) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00100100);
	#1;
	dataIn=12'b110000001001;
	#1;
	if (dataOut==8'b00101001) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00101001);
	#1;
	dataIn=12'b000001000110;
	#1;
	if (dataOut==8'b00110110) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00110110);
	#1;
	dataIn=12'b110101101011;
	#1;
	if (dataOut==8'b00111011) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b00111011);
	#1;
	dataIn=12'b110110011100;
	#1;
	if (dataOut==8'b01000100) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01000100);
	#1;
	dataIn=12'b000010001101;
	#1;
	if (dataOut==8'b01001001) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01001001);
	#1;
	dataIn=12'b110010100100;
	#1;
	if (dataOut==8'b01010110) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01010110);
	#1;
	dataIn=12'b000110111010;
	#1;
	if (dataOut==8'b01011011) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01011011);
	#1;
	dataIn=12'b100011010100;
	#1;
	if (dataOut==8'b01100100) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01100100);
	#1;
	dataIn=12'b010111001001;
	#1;
	if (dataOut==8'b01101001) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01101001);
	#1;
	dataIn=12'b000111100110;
	#1;
	if (dataOut==8'b01110110) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01110110);
	#1;
	dataIn=12'b000011111011;
	#1;
	if (dataOut==8'b01111011) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b01111011);
	#1;
	dataIn=12'b100000010100;
	#1;
	if (dataOut==8'b10000100) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10000100);
	#1;
	dataIn=12'b011100011000;
	#1;
	if (dataOut==8'b10001000) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10001000);
	#1;
	dataIn=12'b101010110111;
	#1;
	if (dataOut==8'b10010111) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10010111);
	#1;
	dataIn=12'b011101101010;
	#1;
	if (dataOut==8'b10011010) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10011010);
	#1;
	dataIn=12'b111001000101;
	#1;
	if (dataOut==8'b10100101) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10100101);
	#1;
	dataIn=12'b001101011000;
	#1;
	if (dataOut==8'b10101000) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10101000);
	#1;
	dataIn=12'b111001100110;
	#1;
	if (dataOut==8'b10110110) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10110110);
	#1;
	dataIn=12'b001101111011;
	#1;
	if (dataOut==8'b10111011) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b10111011);
	#1;
	dataIn=12'b001110010100;
	#1;
	if (dataOut==8'b11000100) result=result+4;
		else $display("time:",$time,":Error in result. For dataIn:%b,  dataOut:%b should be %b",dataIn,dataOut,8'b11000100);


	$display("Result is:%d",result);
	$finish;
	end
endmodule
